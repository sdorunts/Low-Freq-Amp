* C:\Users\sdorunts\Desktop\BMSTU Altium\Low-Freq-Amp\Simulation\Scheme_Sim.sch

* Schematics Version 9.2
* Sat Dec 09 14:44:41 2023


.PARAM         Rn=3 Vhigh=50mV Vlow=-50mV

** Analysis setup **
.tran 0ns 110ms 100ms 10us
.OP 


* From [PSPICE NETLIST] section of C:\Program Files\Orcad\PSpice\PSpice.ini:
.lib "nom.lib"

.INC "Scheme_Sim.net"


.PROBE V(*) I(*) W(*) D(*) NOISE(*) 


.END
